//=====================================================================//
//	Module name: lookup flowKTb in conneciton searcher of UniMon;
//	Communication with lijunnan(lijunnan@nudt.edu.cn)
//	Last edited time: 2018/11/11 (Happy Singles' Day,  Je t'attendrai toujours.)
//	Function outline: UniMan_v1.0
//=====================================================================//

`timescale 1ns/1ps

/**	function description:
*	1) search the flow key table according to the result of hash table;
*		if hiting, return the conneciton table index;
*		otherwise (miss), add a new flow;
*	2) read a free entryID from conf_connTb module (when missing);
*/
module lookup_flowKTb(
reset,
clk,
metadata_in_valid,
metadata_in,
flowK_idx_valid,
flowK_idx_info,
idx_flowKTb,
rdValid_flowKTb,
ctx_flowKTb,
conn_idx_valid,
conn_idx_info,
conn_add_valid,
conn_add_info,
pull_freeFlowID_enable,
free_flowID
);

/*	width or depth or words info of signals
*/
parameter 	w_meta = 113,			// width of metadata, includes hitness(allowTb), flowKey and TCP flag;
			w_key = 104,			// width of flow key;
			w_tcpFlag = 8,			// width of tcp flags, top 2-bit is pad;
			d_connTb = 10,			// depth of connTb;
			w_flowKTb = 120,		// the width of flow key entry, 104b 5-tuple +16b next index;
			d_flowKTb = 10,		// the depth of flow key table;
			d_idxBuffer = 5,			// depth of (flowKTb_conflict) idx buffer, used to buffer meta;
			words_idxBuffer = 32,	// words of idx buffer;
			w_idx = 16,				// width of idx (flowKTb) in idx_flowKIdx_info;
			w_flowID = 16,			// width of flowID;
			w_flowKIdx_info = 16,	// width of flowK_idx_info, i.e., idx_flowKTb;
			w_connIdx_info = 19,	// width of conn_idx_info, include hitness, addness,
									// 	direction, and connection_index ('1' is server2client, '0' is 
									//	client2server);
			w_connAdd_info = 120,	// width of conn_add_info, include flow_key, flowID;

			/* format of 5-tuple in flowKIdx_info, used for comparing with flowKTb */
			b_protocol_key = 96,	// last bit of protocol in flow key;
			b_dstPort_key = 80,		// last bit of dstPort in flow Key;
			b_srcPort_key = 64,		// last bit of srcPort in flow key;
			b_dstIP_key = 32,		// last bit of dstIP in flow key;s
			b_srcIP_key = 0,		// last bit of srcIP in flow key;
			w_proto = 8,			// width of protocol;
			w_ip = 32,				// width of ip;
			w_port = 16,			// width of port;

			b_flowK_flowKTb = 16,	// last bit of the idx_info in flowKTb;
			b_nextIdx_flowKTb = 0,	// last bit of the idx_info in flowKTb;

			SYN_ACK = 8'h12,		// ack & syn;
			ONLY_SYN = 8'h02;		// tcp flag: syn;

input								clk;
input								reset;
input								metadata_in_valid;
input		[w_meta-1:0]			metadata_in;
input								flowK_idx_valid;
input		[w_flowKIdx_info-1:0]	flowK_idx_info;
output	reg	[d_flowKTb-1:0]		idx_flowKTb;
output	reg							rdValid_flowKTb;
input		[w_flowKTb-1:0]		ctx_flowKTb;
output	reg							conn_idx_valid;
output	reg	[w_connIdx_info-1:0]	conn_idx_info;
output	reg							conn_add_valid;
output	reg	[w_connAdd_info-1:0]	conn_add_info;
output	reg							pull_freeFlowID_enable;
input		[w_flowID-1:0]			free_flowID;

/*************************************************************************************/
/***varialbe declaration */
/**	flowKIdx_info buffer */
reg									rdreq_meta;
wire								empty_meta;
wire		[w_meta-1:0]			ctx_meta;

/**	flowKIdx_info buffer */
reg									rdreq_flowKIdx_info;
wire								empty_flowKIdx_info;
wire		[w_flowKIdx_info-1:0]	ctx_flowKIdx_info;

/**	temps used to maintain internal variables
*	flowKey_temp[0] used to save the origirnal 5-tuple info.;
*	flowKey_temp[1] used to save the opposite 5-tuple info.;
*/
reg			[w_key-1:0]				flowKey_temp[1:0];
reg			[w_tcpFlag-1:0]			tcpFlag_temp;
reg									hit_temp;

/**	variables generated by searchFlowKTb;
*	pad_flowID is the difference between the w_flowID and d_flowKTb;
*/
reg 			[w_flowID-1-d_flowKTb:0]	pad_flowID;

/*************************************************************************************/
/***	state register declaration
*/
reg	[3:0]	state_searchFlowKTb;
parameter	IDLE_S				= 4'd0,
			READ_BUFFER_S	= 4'd1,
			WAIT_RAM_1_S		= 4'd2,
			WAIT_RAM_2_S		= 4'd3,
			READ_FLOWKTB_S	= 4'd4,
			ADD_A_FLOW_S	= 4'd5;

/*************************************************************************************/
/***	submodule declaration */
/**	meta_buffer used to cache metadata_in;
*/
fifo_113_32 meta_buffer (
  .clk(clk),      				// input wire clk
  .srst(!reset),    				// input wire srst
  .din(metadata_in),      	// input wire [119 : 0] din
  .wr_en(metadata_in_valid),  // input wire wr_en
  .rd_en(rdreq_meta),  	// input wire rd_en
  .dout(ctx_meta),   		 // output wire [119 : 0] dout
  .full(),    					// output wire full
  .empty(empty_meta)  	// output wire empty
);

/**	flowKIdx_info_buffer used to cache flowK_idx_info;
*/
fifo_16_32 flowKIdx_info_buffer (
  .clk(clk),      						// input wire clk
  .srst(!reset),    						// input wire srst
  .din(flowK_idx_info),      			// input wire [119 : 0] din
  .wr_en(flowK_idx_valid),  			// input wire wr_en
  .rd_en(rdreq_flowKIdx_info),  		// input wire rd_en
  .dout(ctx_flowKIdx_info),   		 // output wire [119 : 0] dout
  .full(),    							// output wire full
  .empty(empty_flowKIdx_info)  	// output wire empty
);
		
/*************************************************************************************/
/**	this state machine is used to search flowKTb;

*	Super day for bench press!
*	If this code has not been updated for a long time, there are two possibilities:
*		1) I was crushed by the barbell;
*		2) The barbell crushed me.
*
*/
always @(posedge clk or negedge reset) begin
	if (!reset) begin
		rdreq_flowKIdx_info <= 1'b0;
		rdreq_meta <= 1'b0;
		conn_add_valid <= 1'b0;
		conn_add_info <= {w_connAdd_info{1'b0}};
		conn_idx_valid <= 1'b0;
		conn_idx_info <= {w_connIdx_info{1'b0}};
		rdValid_flowKTb <= 1'b0;
		idx_flowKTb <= {d_flowKTb{1'b0}};
		pull_freeFlowID_enable <= 1'b0;
		
		state_searchFlowKTb <= IDLE_S;
	end
	else begin
		case(state_searchFlowKTb)
			IDLE_S: begin
				conn_add_valid <=  1'b0;
				conn_idx_valid <= 1'b0;
				if(empty_flowKIdx_info == 1'b0) begin
					rdreq_flowKIdx_info <= 1'b1;
					rdreq_meta <= 1'b1;
					state_searchFlowKTb <= READ_BUFFER_S;
				end
				else begin
					state_searchFlowKTb <= IDLE_S;
				end
			end
			READ_BUFFER_S: begin
				rdreq_flowKIdx_info <= 1'b0;
				rdreq_meta <= 1'b0;
				{hit_temp, flowKey_temp[0], tcpFlag_temp} <= ctx_meta;
				{pad_flowID, idx_flowKTb} <= ctx_flowKIdx_info;
				rdValid_flowKTb <= 1'b1;
				state_searchFlowKTb <= WAIT_RAM_1_S;
			end
			WAIT_RAM_1_S: begin
				rdValid_flowKTb <= 1'b0;
				state_searchFlowKTb <= WAIT_RAM_2_S;
				flowKey_temp[1] <= {
					flowKey_temp[0][b_protocol_key+w_proto-1:b_protocol_key], 
					flowKey_temp[0][b_srcPort_key+w_port-1:b_srcPort_key],
					flowKey_temp[0][b_dstPort_key+w_port-1:b_dstPort_key], 
					flowKey_temp[0][b_srcIP_key+w_ip-1:b_srcIP_key], 
					flowKey_temp[0][b_dstIP_key+w_ip-1:b_dstIP_key]};
			end
			WAIT_RAM_2_S: begin
				state_searchFlowKTb <= READ_FLOWKTB_S;
			end
			READ_FLOWKTB_S: begin
				if(idx_flowKTb == {d_flowKTb{1'b0}}) begin
					/** hashTb miss, and from inbound, just adding a new flowKey; */
					if(((tcpFlag_temp&SYN_ACK) == ONLY_SYN) && (hit_temp == 1'b1)) begin
						pull_freeFlowID_enable <= 1'b1;
						state_searchFlowKTb <= ADD_A_FLOW_S;
					end
					else begin /** not a syn packet, just ignore; */
						state_searchFlowKTb <= IDLE_S;
						conn_idx_valid <= 1'b1;
						conn_idx_info <= {w_connIdx_info{1'b0}};
					end
				end
				else begin
					if(flowKey_temp[0] == ctx_flowKTb[b_flowK_flowKTb+w_key-1:
						b_flowK_flowKTb]) 
					begin /** hit,  addness is '0', direction is '0'; */
						conn_idx_valid <= 1'b1;
						conn_idx_info <= {1'b1,1'b0,1'b0,pad_flowID,idx_flowKTb};
						state_searchFlowKTb <= IDLE_S;
					end
					else if(flowKey_temp[1] == ctx_flowKTb[b_flowK_flowKTb+w_key-1:
						b_flowK_flowKTb]) 
					begin /** hit, addness is '0', direction is 1; */
						conn_idx_valid <= 1'b1;
						conn_idx_info <= {1'b1,1'b0,1'b1,pad_flowID,idx_flowKTb};
						state_searchFlowKTb <= IDLE_S;
					end
					else begin /** miss; */
						if(ctx_flowKTb[b_nextIdx_flowKTb+d_flowKTb-1:b_nextIdx_flowKTb] != {w_idx{1'b0}}) 
						begin
							/** lookup the hash chain; */
							idx_flowKTb <= ctx_flowKTb[b_nextIdx_flowKTb+d_flowKTb-1:
								b_nextIdx_flowKTb];
							rdValid_flowKTb <= 1'b1;
							state_searchFlowKTb <= WAIT_RAM_1_S;
						end
						else begin/** addness is '1', direction is '0' */
							if(((tcpFlag_temp&SYN_ACK) == ONLY_SYN) && (hit_temp == 1'b1))begin
								pull_freeFlowID_enable <= 1'b1;
								state_searchFlowKTb <= ADD_A_FLOW_S;
							end
							else begin /** set '0' and ignore packet */
								state_searchFlowKTb <= IDLE_S;
								conn_idx_valid <= 1'b1;
								conn_idx_info <= {w_connIdx_info{1'b0}};
							end
						end
					end
				end
			end
			ADD_A_FLOW_S: begin 
				/** not a pipeline version, flowKey_temp[0] is the 5-tuple */
				pull_freeFlowID_enable <= 1'b0;
				conn_add_valid <= 1'b1;
				conn_add_info <= {flowKey_temp[0],free_flowID};
				conn_idx_valid <= 1'b1;
				conn_idx_info <=  {1'b0,1'b1,1'b0, free_flowID};
				state_searchFlowKTb <= IDLE_S;
			end
			default: begin
				state_searchFlowKTb <= IDLE_S;
			end
		endcase
	end
end

endmodule    
